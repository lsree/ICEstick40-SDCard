`timescale 1ns/1ns

module blinky_tb;
reg clk;
wire LED1, LED2, LED3, LED4, LED5;
wire RLED1, RLED2, RLED3, RLED4, RLED5;

assign {LED1, LED2, LED3, LED4, LED5} = 0;


initial begin
    clk = 0;
end

blinky test_blink(clk, LED1, LED2, LED3, LED4, LED5);
LED_Rotation test_rotation(clk, RLED1, RLED2, RLED3, RLED4, RLED5);

always #1 clk = !clk;

endmodule